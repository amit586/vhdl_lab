`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:07:55 09/23/2020 
// Design Name: 
// Module Name:    fourbitadder 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module fourbitadder(
    input x,
    input y,
    input [3:0] in,
    input carryin,
    output [3:0] sum,
    output carryout
    );


endmodule
